//////////////////////////////////////////////////////////////////////////////
//             Fetching and prepare instruction for execution               //
/////////////////////////////////////////////////////////////////////////////

